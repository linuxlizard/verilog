`define KP_0 8'h70
`define KP_1 8'h71
`define KP_2 8'h72
`define KP_3 8'h73
`define KP_4 8'h74
`define KP_5 8'h75
`define KP_6 8'h76
`define KP_7 8'h77
`define KP_8 8'h78
`define KP_9 8'h79
`define KP_STAR 8'h7c
`define KP_MINUS 8'h7b


