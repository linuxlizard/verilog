`define MUX_SEL_REGISTER_2_LSB 0
`define MUX_SEL_REGISTER_2_MSB 1
`define MUX_SEL_COUNTER_VALUE  2
`define MUX_SEL_COUNTER_CARRY  3
