`define KP_0 8'h70
`define KP_1 8'h69
`define KP_2 8'h72
`define KP_3 8'h7a
`define KP_4 8'h6b
`define KP_5 8'h73
`define KP_6 8'h74
`define KP_7 8'h6c
`define KP_8 8'h75
`define KP_9 8'h7d
`define KP_STAR 8'h7c
`define KP_MINUS 8'h7b

`define KP_KEY_RELEASED 8'hf0

`define KP_0_BCD 4'h0
`define KP_1_BCD 4'h1
`define KP_2_BCD 4'h2
`define KP_3_BCD 4'h3
`define KP_4_BCD 4'h4
`define KP_5_BCD 4'h5
`define KP_6_BCD 4'h6
`define KP_7_BCD 4'h7
`define KP_8_BCD 4'h8
`define KP_9_BCD   4'h9

`define KP_INVALID 8'hff

