`define KP_0 8'h70
`define KP_1 8'h69
`define KP_2 8'h72
`define KP_3 8'h7a
`define KP_4 8'h6b
`define KP_5 8'h73
`define KP_6 8'h74
`define KP_7 8'h6c
`define KP_8 8'h75
`define KP_9 8'h7d
`define KP_STAR 8'h7c
`define KP_MINUS 8'h7b

`define KP_KEY_RELEASED 8'hf0

`define KP_0_BCD 8'h00
`define KP_1_BCD 8'h01
`define KP_2_BCD 8'h02
`define KP_3_BCD 8'h03
`define KP_4_BCD 8'h04
`define KP_5_BCD 8'h05
`define KP_6_BCD 8'h06
`define KP_7_BCD 8'h07
`define KP_8_BCD 8'h08
`define KP_9_BCD   8'h09

//`define KP_STAR_BCD 8'h0a
//`define KP_MINUS_BCD 8'h0b
//`define KP_KEY_RELEASED_BCD 8'hf0

`define KP_INVALID 8'hff

