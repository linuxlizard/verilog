
/* values for PIC readwrite bit */
`define RW_READ 1'b1
`define RW_WRITE 1'b0

/* register values; used with the PIC select bits */
`define SEL_OCR 2'b00
`define SEL_IMR 2'b01
`define SEL_IRR 2'b10
`define SEL_ISR 2'b11
